module user_uart2udp(
    input        clk,            // ϵͳʱ��
    input        rst_n,          // ϵͳ��λ������Ч
    
    input        uart_rx_done,   // UART��������ź�
    input [7:0]  uart_rx_data,   // UART���յ�������

    output reg   rec_en,         // ����ʹ���ź�
    output reg [7:0] rec_data,   // ���յ�������
    output reg   tx_start_en     // UDP���������ź�
);

always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        rec_en       <= 1'b0;
        rec_data     <= 8'b0;
        tx_start_en  <= 1'b0;
    end else begin
        rec_en       <= uart_rx_done;          // �����յ�����ʱ��ʹ�ܽ����ź�
        rec_data     <= uart_rx_data;          // �洢���յ�������

        if (uart_rx_done && (uart_rx_data == 8'h0A)) begin  // ����յ����з�������UDP����
            tx_start_en <= 1'b1;
        end else begin
            tx_start_en <= 1'b0;
        end
    end
end

endmodule